[HTMLEFS][1][Asana Client][Enterprise, VMC , Test][Asana Client; Created by Derry Everson 04/10/2020][Asana Client][//localserver/EncounterForms/HtmlForms/Asana-Client/index.html][Arial]
